// -------------------------------------------------------
// -- StageRegWB.v - Stage register of WB
// -------------------------------------------------------
// Bugen Zhao 2020
// -------------------------------------------------------

`timescale 1ns / 1ps
`include "ISA.v"

module StageRegWB(
           input clk,

           input wire [`WORD] memNewPC, memInstruction,
           input wire [`WORD] memAluOut, memMemOut,
           input wire [ `REG] memWriteReg,
           input wire         memMemRead,

           output reg [`WORD] wbNewPC, wbInstruction,
           output reg [`WORD] wbAluOut, wbMemOut,
           output reg [ `REG] wbWriteReg,
           output reg         wbMemRead
       );

// reg [`WORD] newPC, instruction;
// reg [`WORD] aluOut, memOut;
// reg [ `REG] writeReg;
// reg         memRead;

always @(negedge clk) begin
    wbNewPC = memNewPC;
    wbInstruction = memInstruction;
    wbAluOut = memAluOut;
    wbMemOut = memMemOut;
    wbWriteReg = memWriteReg;
    wbMemRead = memMemRead;
end

// assign wbNewPC = newPC;
// assign wbInstruction = instruction;
// assign wbAluOut = aluOut;
// assign wbMemOut = memOut;
// assign wbWriteReg = writeReg;
// assign wbMemRead = memRead;

endmodule // StageRegWB
